module main(sw0 , led0, led);

input sw0;
output led0;
output reg [7:0] led;

assign led0 = sw0;



endmodule

